module calculadora_sincrona(
    input [7:0] entrada,
    input [2:0] codigo,
    output reg [7:0] saida
);
    
//insira seu código aqui

endmodule